interface uart_if(

    input logic clk
);
    logic rx;
    logic tx;

endinterface