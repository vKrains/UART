package uvm_uart_test_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "../uvma_apb/dv/uvma_apb/src/uvma_apb_plg.sv"
    `include "../../src/AXIS_UVM_Agent/src/axis_intf.sv"
    `include "../../src/AXIS_UVM_Agent/src/axis_include.svh"
    `include "uvm_uart_env.sv"
    `include "uvm_uart_base_test.sv"
    
endpackage