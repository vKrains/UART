class uart_sequence_item extends uvm_sequence_item;
  `uvm_object_utils(uart_sequence_item)


endclass
